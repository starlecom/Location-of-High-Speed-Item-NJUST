library verilog;
use verilog.vl_types.all;
entity topdesign_vlg_vec_tst is
end topdesign_vlg_vec_tst;
